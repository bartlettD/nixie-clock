** Profile: "Basic Flyback-TPS40210"  [ c:\users\dylan\nixie-clock\simulation\flyback\flyback-PSpiceFiles\Basic Flyback\TPS40210.sim ] 

** Creating circuit file "TPS40210.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../SBR1U400P1.spice.lib" 
.LIB "../../../p_se50paj.lib" 
.LIB "../../../dmt6030lfcl.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS THREADS= 1
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\Basic Flyback.net" 


.END
