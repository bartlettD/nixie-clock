** Profile: "TPS55330-TPS55330-tran"  [ C:\Users\dylan\nixie-clock\Simulation\flyback\flyback-pspicefiles\tps55330\tps55330-tran.sim ] 

** Creating circuit file "TPS55330-tran.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS ABSTOL= 10n
.OPTIONS ITL1= 1500
.OPTIONS ITL2= 400
.OPTIONS ITL4= 400
.OPTIONS VNTOL= 10u
.OPTIONS THREADS= 1
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\TPS55330.net" 


.END
