** Profile: "LM5155-lm5155"  [ c:\users\dylan\nixie-clock\simulation\flyback\flyback-pspicefiles\lm5155\lm5155.sim ] 

** Creating circuit file "lm5155.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../WE-FLYLT.lib" 
.LIB "../../../SBR1U400P1.spice.lib" 
.LIB "../../../p_se50paj.lib" 
.LIB "../../../dmt6030lfcl.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5m 0 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.PROBE64 N([N27760])
.PROBE64 N([N28164])
.PROBE64 I(L_L1)
.INC "..\LM5155.net" 


.END
