** Profile: "Basic Flyback-transient"  [ C:\Users\dylan\nixie-clock\Simulation\flyback\flyback-pspicefiles\basic flyback\transient.sim ] 

** Creating circuit file "transient.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../dmt6030lfcl.lib" 
* From [PSPICE NETLIST] section of C:\cds_spb_home\cdssetup\OrCAD_PSpiceTIPSpice_Install\23.1.0\PSpice.ini file:
.lib "nom_pspti.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 30m 0 
.OPTIONS ADVCONV
.OPTIONS FILEMODELSEARCH
.OPTIONS THREADS= 1
.PROBE64 N([N14510])
.PROBE64 W(X_U1)
.PROBE64 N([N14585])
.INC "..\Basic Flyback.net" 


.END
